module cpu_tb
endmodule